library verilog;
use verilog.vl_types.all;
entity sim is
end sim;
